module register(src0, src1, dst, we, data, clk, rst_n, outa, outb);
	input clk, rst_n;
	input [5:0] dst;
	input we;
	input [44:0] data;
  input [5:0] src0, src1;
	output [44:0] outa, outb;

	wire [44:0] MONDAI, KOTAE;

	reg [44:0] regis [61:0];
  reg [44:0] answer;
	parameter [44:0] BOARD0 = 45'b000000000000000000000000000_000_001_010_011_100_101,
    BOARD1 = 45'b000000000000000000000000000_000_001_011_100_010_101,
    BOARD2 = 45'b000000000000000000000000000_000_001_100_010_011_101,
    BOARD3 = 45'b000000000000000000000000000_000_010_001_100_011_101,
    BOARD4 = 45'b000000000000000000000000000_000_010_011_001_100_101,
    BOARD5 = 45'b000000000000000000000000000_000_010_100_011_001_101,
    BOARD6 = 45'b000000000000000000000000000_000_011_001_010_100_101,
    BOARD7 = 45'b000000000000000000000000000_000_011_010_100_001_101,
    BOARD8 = 45'b000000000000000000000000000_000_011_100_001_010_101,
    BOARD9 = 45'b000000000000000000000000000_000_100_001_011_010_101,
    BOARD10 = 45'b000000000000000000000000000_000_100_010_001_011_101,
    BOARD11 = 45'b000000000000000000000000000_000_100_011_010_001_101,
    BOARD12 = 45'b000000000000000000000000000_001_000_010_100_011_101,
    BOARD13 = 45'b000000000000000000000000000_001_000_011_010_100_101,
    BOARD14 = 45'b000000000000000000000000000_001_000_100_011_010_101,
    BOARD15 = 45'b000000000000000000000000000_001_010_000_011_100_101,
    BOARD16 = 45'b000000000000000000000000000_001_010_011_100_000_101,
    BOARD17 = 45'b000000000000000000000000000_001_010_100_000_011_101,
    BOARD18 = 45'b000000000000000000000000000_001_011_000_100_010_101,
    BOARD19 = 45'b000000000000000000000000000_001_011_010_000_100_101,
    BOARD20 = 45'b000000000000000000000000000_001_011_100_010_000_101,
    BOARD21 = 45'b000000000000000000000000000_001_100_000_010_011_101,
    BOARD22 = 45'b000000000000000000000000000_001_100_010_011_000_101,
    BOARD23 = 45'b000000000000000000000000000_001_100_011_000_010_101,
    BOARD24 = 45'b000000000000000000000000000_010_000_001_011_100_101,
    BOARD25 = 45'b000000000000000000000000000_010_000_011_100_001_101,
    BOARD26 = 45'b000000000000000000000000000_010_000_100_001_011_101,
    BOARD27 = 45'b000000000000000000000000000_010_001_000_100_011_101,
    BOARD28 = 45'b000000000000000000000000000_010_001_011_000_100_101,
    BOARD29 = 45'b000000000000000000000000000_010_001_100_011_000_101,
    BOARD30 = 45'b000000000000000000000000000_010_011_000_001_100_101,
    BOARD31 = 45'b000000000000000000000000000_010_011_001_100_000_101,
    BOARD32 = 45'b000000000000000000000000000_010_011_100_000_001_101,
    BOARD33 = 45'b000000000000000000000000000_010_100_000_011_001_101,
    BOARD34 = 45'b000000000000000000000000000_010_100_001_000_011_101,
    BOARD35 = 45'b000000000000000000000000000_010_100_011_001_000_101,
    BOARD36 = 45'b000000000000000000000000000_011_000_001_100_010_101,
    BOARD37 = 45'b000000000000000000000000000_011_000_010_001_100_101,
    BOARD38 = 45'b000000000000000000000000000_011_000_100_010_001_101,
    BOARD39 = 45'b000000000000000000000000000_011_001_000_010_100_101,
    BOARD40 = 45'b000000000000000000000000000_011_001_010_100_000_101,
    BOARD41 = 45'b000000000000000000000000000_011_001_100_000_010_101,
    BOARD42 = 45'b000000000000000000000000000_011_010_000_100_001_101,
    BOARD43 = 45'b000000000000000000000000000_011_010_001_000_100_101,
    BOARD44 = 45'b000000000000000000000000000_011_010_100_001_000_101,
    BOARD45 = 45'b000000000000000000000000000_011_100_000_001_010_101,
    BOARD46 = 45'b000000000000000000000000000_011_100_001_010_000_101,
    BOARD47 = 45'b000000000000000000000000000_011_100_010_000_001_101,
    BOARD48 = 45'b000000000000000000000000000_100_000_001_010_011_101,
    BOARD49 = 45'b000000000000000000000000000_100_000_010_011_001_101,
    BOARD50 = 45'b000000000000000000000000000_100_000_011_001_010_101,
    BOARD51 = 45'b000000000000000000000000000_100_001_000_011_010_101,
    BOARD52 = 45'b000000000000000000000000000_100_001_010_000_011_101,
    BOARD53 = 45'b000000000000000000000000000_100_001_011_010_000_101,
    BOARD54 = 45'b000000000000000000000000000_100_010_000_001_011_101,
    BOARD55 = 45'b000000000000000000000000000_100_010_001_011_000_101,
    BOARD56 = 45'b000000000000000000000000000_100_010_011_000_001_101,
    BOARD57 = 45'b000000000000000000000000000_100_011_000_010_001_101,
    BOARD58 = 45'b000000000000000000000000000_100_011_001_000_010_101,
    BOARD59 = 45'b000000000000000000000000000_100_011_010_001_000_101,
    QUESTION = 45'b000000000000000000000000000_000_001_011_100_010_101;
	
	always @(posedge clk) begin
		if (!rst_n) begin
			// $B=i4|!&8=:_$NHWLL(B
			// ####_1111_2222_3333_4444_5555_7777
			regis[0] <= BOARD0;
			regis[1] <= BOARD1;
			regis[2] <= BOARD2;
			regis[3] <= BOARD3;
			regis[4] <= BOARD4;
			regis[5] <= BOARD5;
			regis[6] <= BOARD6;
			regis[7] <= BOARD7;
			regis[8] <= BOARD8;
			regis[9] <= BOARD9;
			regis[10] <= BOARD10;
			regis[11] <= BOARD11;
			regis[12] <= BOARD12;
			regis[13] <= BOARD13;
			regis[14] <= BOARD14;
			regis[15] <= BOARD15;
			regis[16] <= BOARD16;
			regis[17] <= BOARD17;
			regis[18] <= BOARD18;
			regis[19] <= BOARD19;
			regis[20] <= BOARD20;
			regis[21] <= BOARD21;
			regis[22] <= BOARD22;
			regis[23] <= BOARD23;
			regis[24] <= BOARD24;
			regis[25] <= BOARD25;
			regis[26] <= BOARD26;
			regis[27] <= BOARD27;
			regis[28] <= BOARD28;
			regis[29] <= BOARD29;
			regis[30] <= BOARD30;
			regis[31] <= BOARD31;
			regis[32] <= BOARD32;
			regis[33] <= BOARD33;
			regis[34] <= BOARD34;
			regis[35] <= BOARD35;
			regis[36] <= BOARD36;
			regis[37] <= BOARD37;
			regis[38] <= BOARD38;
			regis[39] <= BOARD39;
			regis[40] <= BOARD40;
			regis[41] <= BOARD41;
			regis[42] <= BOARD42;
			regis[43] <= BOARD43;
			regis[44] <= BOARD44;
			regis[45] <= BOARD45;
			regis[46] <= BOARD46;
			regis[47] <= BOARD47;
			regis[48] <= BOARD48;
			regis[49] <= BOARD49;
			regis[50] <= BOARD50;
			regis[51] <= BOARD51;
			regis[52] <= BOARD52;
			regis[53] <= BOARD53;
			regis[54] <= BOARD54;
			regis[55] <= BOARD55;
			regis[56] <= BOARD56;
			regis[57] <= BOARD57;
			regis[58] <= BOARD58;
			regis[59] <= BOARD59;
      regis[60] <= QUESTION;
      regis[61] <= 0;
		end else begin
			if (we) begin
				regis[dst] <= data;
			end else begin
				regis[dst] <= regis[dst];
			end
		end
	end

	assign outa = regis[src0];
	assign outb = regis[src1];
	assign MONDAI = regis[60];
	assign KOTAE = regis[61];
endmodule
